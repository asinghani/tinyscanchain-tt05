`default_nettype none

module tt_um_asinghani_tinyscanchain_tt05 (
    input  wire [7:0] ui_in,    // Dedicated inputs - connected to the input switches
    output wire [7:0] uo_out,   // Dedicated outputs - connected to the 7 segment display
    input  wire [7:0] uio_in,   // IOs: Bidirectional Input path
    output wire [7:0] uio_out,  // IOs: Bidirectional Output path
    output wire [7:0] uio_oe,   // IOs: Bidirectional Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // will go high when the design is enabled
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

    seven_segment_seconds mod (
        .clk(clk),
        .rst(!rst_n),
        .ena(ui_in[0]),
        .led_out(uo_out[6:0]),
        
        .scan_in(ui_in[1]),
        .scan_en(ui_in[2]),
        .scan_out(uo_out[7])
    );

    assign uio_out = '0;
    assign uio_oe  = '0;

endmodule
